module RAM #(parameter USER_CAPACITY, parameter ASSET_COUNT)(
    input wire [15:0] name,
    input wire 
)
parameter LOG = $clog(USER_CAPACITY);


endmodule

module RAM_Instruction_fetch